// nios.v

// Generated using ACDS version 17.0 602

`timescale 1 ps / 1 ps
module nios (
		input  wire       clk_clk,                        //                        clk.clk
		output wire [7:0] led_external_connection_export, //    led_external_connection.export
		input  wire       reset_reset_n,                  //                      reset.reset_n
		input  wire       uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire       uart_0_external_connection_txd  //                           .txd
	);

	wire         nios2_gen2_0_custom_instruction_master_readra;                                   // nios2_gen2_0:D_ci_readra -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_a;                                        // nios2_gen2_0:D_ci_a -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_b;                                        // nios2_gen2_0:D_ci_b -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_gen2_0_custom_instruction_master_c;                                        // nios2_gen2_0:D_ci_c -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_readrb;                                   // nios2_gen2_0:D_ci_readrb -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_readrb
	wire         nios2_gen2_0_custom_instruction_master_clk;                                      // nios2_gen2_0:E_ci_multi_clock -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_gen2_0_custom_instruction_master_ipending;                                 // nios2_gen2_0:W_ci_ipending -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_ipending
	wire         nios2_gen2_0_custom_instruction_master_start;                                    // nios2_gen2_0:E_ci_multi_start -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios2_gen2_0_custom_instruction_master_reset_req;                                // nios2_gen2_0:E_ci_multi_reset_req -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_gen2_0_custom_instruction_master_done;                                     // nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_done -> nios2_gen2_0:E_ci_multi_done
	wire   [7:0] nios2_gen2_0_custom_instruction_master_n;                                        // nios2_gen2_0:D_ci_n -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_result;                                   // nios2_gen2_0_custom_instruction_master_translator:ci_slave_result -> nios2_gen2_0:E_ci_result
	wire         nios2_gen2_0_custom_instruction_master_estatus;                                  // nios2_gen2_0:W_ci_estatus -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_estatus
	wire         nios2_gen2_0_custom_instruction_master_clk_en;                                   // nios2_gen2_0:E_ci_multi_clk_en -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] nios2_gen2_0_custom_instruction_master_datab;                                    // nios2_gen2_0:E_ci_datab -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_dataa;                                    // nios2_gen2_0:E_ci_dataa -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_reset;                                    // nios2_gen2_0:E_ci_multi_reset -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_gen2_0_custom_instruction_master_writerc;                                  // nios2_gen2_0:D_ci_writerc -> nios2_gen2_0_custom_instruction_master_translator:ci_slave_writerc
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra;        // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readra -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a;             // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_a -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b;             // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_b -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk;           // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clk -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb;        // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c;             // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_c -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_start -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n;             // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_n -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_clken -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_datab -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset;         // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_reset -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc;       // nios2_gen2_0_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result; // div_0:result -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_clk -> div_0:clk
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_clken -> div_0:clk_en
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_datab -> div_0:datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> div_0:dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_start -> div_0:start
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_reset -> div_0:reset
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done;   // div_0:done -> nios2_gen2_0_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readra;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_readra -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_a;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_a -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_b;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_b -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_readrb -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_c;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_c -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk;            // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_clk -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending;       // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_ipending -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_start;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_start -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req;      // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_done;           // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_done -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_n;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_n -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_result;         // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_result -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_estatus -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_clken -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_datab;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_datab -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_dataa -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_reset -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master1_writerc -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_result; // mult_0:result -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk;    // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_clk -> mult_0:clk
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en; // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_clken -> mult_0:clk_en
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_datab -> mult_0:datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> mult_0:dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_start;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_start -> mult_0:start
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_reset -> mult_0:reset
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_done;   // mult_0:done -> nios2_gen2_0_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readra;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_readra -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_readra
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_a;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_a -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_a
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_b;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_b -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_b
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readrb;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_readrb -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_readrb
	wire   [4:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_c;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_c -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_c
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk;            // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_clk -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_clk
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_ipending;       // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_ipending -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_ipending
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_start;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_start -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_start
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset_req;      // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_reset_req -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_reset_req
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_done;           // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_done -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_done
	wire   [7:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_n;              // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_n -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_n
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_result;         // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_result -> nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_result
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_estatus;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_estatus -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_estatus
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk_en;         // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_clken -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_clken
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_datab;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_datab -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_dataa;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_dataa -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset;          // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_reset -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_reset
	wire         nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_writerc;        // nios2_gen2_0_custom_instruction_master_multi_xconnect:ci_master2_writerc -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_slave_writerc
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_result; // resto_0:result -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_result
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk;    // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_clk -> resto_0:clk
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk_en; // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_clken -> resto_0:clk_en
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_datab;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_datab -> resto_0:datab
	wire  [31:0] nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_dataa;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_dataa -> resto_0:dataa
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_start;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_start -> resto_0:start
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_reset;  // nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_reset -> resto_0:reset
	wire         nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_done;   // resto_0:done -> nios2_gen2_0_custom_instruction_master_multi_slave_translator2:ci_master_done
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                               // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                            // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                            // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [13:0] nios2_gen2_0_data_master_address;                                                // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                             // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                   // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                                  // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                              // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                        // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                     // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [13:0] nios2_gen2_0_instruction_master_address;                                         // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                            // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                         // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                      // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_uart_0_s1_chipselect;                                          // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                                            // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                                             // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_read;                                                // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                                       // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire         mm_interconnect_0_uart_0_s1_write;                                               // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                                           // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire         mm_interconnect_0_led_s1_chipselect;                                             // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                               // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                                // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                                  // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                              // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                  // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                   // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                     // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                 // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                     // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                                        // uart_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                            // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                                  // rst_controller:reset_out -> [irq_mapper:reset, led:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, uart_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                              // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                                          // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1

	div div_0 (
		.dataa  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                              .datab
		.result (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.clk    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                              .clk
		.clk_en (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.start  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.reset  (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.done   (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done)    //                              .done
	);

	nios_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	mul mult_0 (
		.dataa  (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab  (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                              .datab
		.result (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_result), //                              .result
		.clk    (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //                              .clk
		.clk_en (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //                              .clk_en
		.start  (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                              .start
		.reset  (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //                              .reset
		.done   (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_done)    //                              .done
	);

	nios_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (nios2_gen2_0_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (nios2_gen2_0_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (nios2_gen2_0_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (nios2_gen2_0_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (nios2_gen2_0_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_gen2_0_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_gen2_0_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_gen2_0_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_gen2_0_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_gen2_0_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_gen2_0_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_gen2_0_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_gen2_0_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (nios2_gen2_0_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (nios2_gen2_0_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (nios2_gen2_0_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (nios2_gen2_0_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_gen2_0_custom_instruction_master_ipending)             //                          .ipending
	);

	nios_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	resto resto_0 (
		.dataa  (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab  (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_datab),  //                              .datab
		.result (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_result), //                              .result
		.clk    (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk),    //                              .clk
		.clk_en (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk_en), //                              .clk_en
		.start  (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_start),  //                              .start
		.reset  (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_reset),  //                              .reset
		.done   (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_done)    //                              .done
	);

	nios_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),            // external_connection.export
		.txd           (uart_0_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver0_irq)                   //                 irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_gen2_0_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_gen2_0_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_gen2_0_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_gen2_0_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_gen2_0_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_gen2_0_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_gen2_0_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_gen2_0_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_gen2_0_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_gen2_0_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_gen2_0_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_gen2_0_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_gen2_0_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_gen2_0_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_gen2_0_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_gen2_0_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_gen2_0_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_gen2_0_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_gen2_0_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                            //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                            //                .datab
		.comb_ci_master_result     (),                                                                            //                .result
		.comb_ci_master_n          (),                                                                            //                .n
		.comb_ci_master_readra     (),                                                                            //                .readra
		.comb_ci_master_readrb     (),                                                                            //                .readrb
		.comb_ci_master_writerc    (),                                                                            //                .writerc
		.comb_ci_master_a          (),                                                                            //                .a
		.comb_ci_master_b          (),                                                                            //                .b
		.comb_ci_master_c          (),                                                                            //                .c
		.comb_ci_master_ipending   (),                                                                            //                .ipending
		.comb_ci_master_estatus    (),                                                                            //                .estatus
		.multi_ci_master_clk       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                        //     (terminated)
		.ci_slave_multi_result     (),                                                                            //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                                 //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                        //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                    //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                    //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                                     //     (terminated)
	);

	nios_nios2_gen2_0_custom_instruction_master_multi_xconnect nios2_gen2_0_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                            //           .ipending
		.ci_slave_estatus     (),                                                                            //           .estatus
		.ci_slave_clk         (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_gen2_0_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_done),       //           .done
		.ci_master2_dataa     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_dataa),      // ci_master2.dataa
		.ci_master2_datab     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_datab),      //           .datab
		.ci_master2_result    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_result),     //           .result
		.ci_master2_n         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_n),          //           .n
		.ci_master2_readra    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readra),     //           .readra
		.ci_master2_readrb    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readrb),     //           .readrb
		.ci_master2_writerc   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_writerc),    //           .writerc
		.ci_master2_a         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_a),          //           .a
		.ci_master2_b         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_b),          //           .b
		.ci_master2_c         (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_c),          //           .c
		.ci_master2_ipending  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_ipending),   //           .ipending
		.ci_master2_estatus   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_estatus),    //           .estatus
		.ci_master2_clk       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk),        //           .clk
		.ci_master2_reset     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset),      //           .reset
		.ci_master2_clken     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk_en),     //           .clk_en
		.ci_master2_reset_req (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset_req),  //           .reset_req
		.ci_master2_start     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_start),      //           .start
		.ci_master2_done      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_0_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_gen2_0_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                                // (terminated)
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   (),                                                                                // (terminated)
		.ci_master_reset_req ()                                                                                 // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_0_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios2_gen2_0_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_n         (),                                                                                // (terminated)
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   (),                                                                                // (terminated)
		.ci_master_reset_req ()                                                                                 // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_gen2_0_custom_instruction_master_multi_slave_translator2 (
		.ci_slave_dataa      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_datab),          //          .datab
		.ci_slave_result     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_result),         //          .result
		.ci_slave_n          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_n),              //          .n
		.ci_slave_readra     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readra),         //          .readra
		.ci_slave_readrb     (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_writerc),        //          .writerc
		.ci_slave_a          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_a),              //          .a
		.ci_slave_b          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_b),              //          .b
		.ci_slave_c          (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_c),              //          .c
		.ci_slave_ipending   (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_estatus),        //          .estatus
		.ci_slave_clk        (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk),            //          .clk
		.ci_slave_clken      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_reset),          //          .reset
		.ci_slave_start      (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_start),          //          .start
		.ci_slave_done       (nios2_gen2_0_custom_instruction_master_multi_xconnect_ci_master2_done),           //          .done
		.ci_master_dataa     (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_result), //          .result
		.ci_master_clk       (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_start),  //          .start
		.ci_master_done      (nios2_gen2_0_custom_instruction_master_multi_slave_translator2_ci_master_done),   //          .done
		.ci_master_n         (),                                                                                // (terminated)
		.ci_master_readra    (),                                                                                // (terminated)
		.ci_master_readrb    (),                                                                                // (terminated)
		.ci_master_writerc   (),                                                                                // (terminated)
		.ci_master_a         (),                                                                                // (terminated)
		.ci_master_b         (),                                                                                // (terminated)
		.ci_master_c         (),                                                                                // (terminated)
		.ci_master_ipending  (),                                                                                // (terminated)
		.ci_master_estatus   (),                                                                                // (terminated)
		.ci_master_reset_req ()                                                                                 // (terminated)
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                    //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                           //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                       //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                        //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                              //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                          //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                             //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                         //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                       //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                    //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                       //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                   //                                         .readdata
		.led_s1_address                                 (mm_interconnect_0_led_s1_address),                           //                                   led_s1.address
		.led_s1_write                                   (mm_interconnect_0_led_s1_write),                             //                                         .write
		.led_s1_readdata                                (mm_interconnect_0_led_s1_readdata),                          //                                         .readdata
		.led_s1_writedata                               (mm_interconnect_0_led_s1_writedata),                         //                                         .writedata
		.led_s1_chipselect                              (mm_interconnect_0_led_s1_chipselect),                        //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                                         .debugaccess
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),              //                      onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                //                                         .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),             //                                         .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),            //                                         .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),           //                                         .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),           //                                         .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                //                                         .clken
		.uart_0_s1_address                              (mm_interconnect_0_uart_0_s1_address),                        //                                uart_0_s1.address
		.uart_0_s1_write                                (mm_interconnect_0_uart_0_s1_write),                          //                                         .write
		.uart_0_s1_read                                 (mm_interconnect_0_uart_0_s1_read),                           //                                         .read
		.uart_0_s1_readdata                             (mm_interconnect_0_uart_0_s1_readdata),                       //                                         .readdata
		.uart_0_s1_writedata                            (mm_interconnect_0_uart_0_s1_writedata),                      //                                         .writedata
		.uart_0_s1_begintransfer                        (mm_interconnect_0_uart_0_s1_begintransfer),                  //                                         .begintransfer
		.uart_0_s1_chipselect                           (mm_interconnect_0_uart_0_s1_chipselect)                      //                                         .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
