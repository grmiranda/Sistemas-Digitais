// proj_qsys.v

// Generated using ACDS version 13.1 182 at 2019.04.08.22:31:22

`timescale 1 ps / 1 ps
module proj_qsys (
		input  wire       clk_clk,                            //                         clk.clk
		input  wire [3:0] buttons_external_connection_export, // buttons_external_connection.export
		output wire [3:0] leds_external_connection_export,    //    leds_external_connection.export
		output wire       en_export,                          //                          en.export
		output wire       rw_export,                          //                          rw.export
		output wire       rs_export,                          //                          rs.export
		output wire [7:0] db_export                           //                          db.export
	);

	wire         nios_jtag_debug_module_reset_reset;                                      // nios:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	wire  [31:0] nios_custom_instruction_master_result;                                   // nios_custom_instruction_master_translator:ci_slave_result -> nios:E_ci_result
	wire   [4:0] nios_custom_instruction_master_b;                                        // nios:D_ci_b -> nios_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_c;                                        // nios:D_ci_c -> nios_custom_instruction_master_translator:ci_slave_c
	wire         nios_custom_instruction_master_done;                                     // nios_custom_instruction_master_translator:ci_slave_multi_done -> nios:E_ci_multi_done
	wire         nios_custom_instruction_master_clk_en;                                   // nios:E_ci_multi_clk_en -> nios_custom_instruction_master_translator:ci_slave_multi_clken
	wire   [4:0] nios_custom_instruction_master_a;                                        // nios:D_ci_a -> nios_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_n;                                        // nios:D_ci_n -> nios_custom_instruction_master_translator:ci_slave_n
	wire         nios_custom_instruction_master_writerc;                                  // nios:D_ci_writerc -> nios_custom_instruction_master_translator:ci_slave_writerc
	wire         nios_custom_instruction_master_clk;                                      // nios:E_ci_multi_clock -> nios_custom_instruction_master_translator:ci_slave_multi_clk
	wire         nios_custom_instruction_master_reset_req;                                // nios:E_ci_multi_reset_req -> nios_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios_custom_instruction_master_start;                                    // nios:E_ci_multi_start -> nios_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] nios_custom_instruction_master_dataa;                                    // nios:E_ci_dataa -> nios_custom_instruction_master_translator:ci_slave_dataa
	wire         nios_custom_instruction_master_readra;                                   // nios:D_ci_readra -> nios_custom_instruction_master_translator:ci_slave_readra
	wire         nios_custom_instruction_master_reset;                                    // nios:E_ci_multi_reset -> nios_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] nios_custom_instruction_master_datab;                                    // nios:E_ci_datab -> nios_custom_instruction_master_translator:ci_slave_datab
	wire         nios_custom_instruction_master_readrb;                                   // nios:D_ci_readrb -> nios_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_result;        // nios_custom_instruction_master_multi_xconnect:ci_slave_result -> nios_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_b;             // nios_custom_instruction_master_translator:multi_ci_master_b -> nios_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_c;             // nios_custom_instruction_master_translator:multi_ci_master_c -> nios_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] nios_custom_instruction_master_translator_multi_ci_master_a;             // nios_custom_instruction_master_translator:multi_ci_master_a -> nios_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk_en;        // nios_custom_instruction_master_translator:multi_ci_master_clken -> nios_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         nios_custom_instruction_master_translator_multi_ci_master_done;          // nios_custom_instruction_master_multi_xconnect:ci_slave_done -> nios_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios_custom_instruction_master_translator_multi_ci_master_n;             // nios_custom_instruction_master_translator:multi_ci_master_n -> nios_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         nios_custom_instruction_master_translator_multi_ci_master_writerc;       // nios_custom_instruction_master_translator:multi_ci_master_writerc -> nios_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios_custom_instruction_master_translator_multi_ci_master_clk;           // nios_custom_instruction_master_translator:multi_ci_master_clk -> nios_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset_req;     // nios_custom_instruction_master_translator:multi_ci_master_reset_req -> nios_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios_custom_instruction_master_translator_multi_ci_master_start;         // nios_custom_instruction_master_translator:multi_ci_master_start -> nios_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_dataa;         // nios_custom_instruction_master_translator:multi_ci_master_dataa -> nios_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios_custom_instruction_master_translator_multi_ci_master_readra;        // nios_custom_instruction_master_translator:multi_ci_master_readra -> nios_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         nios_custom_instruction_master_translator_multi_ci_master_reset;         // nios_custom_instruction_master_translator:multi_ci_master_reset -> nios_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_translator_multi_ci_master_datab;         // nios_custom_instruction_master_translator:multi_ci_master_datab -> nios_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         nios_custom_instruction_master_translator_multi_ci_master_readrb;        // nios_custom_instruction_master_translator:multi_ci_master_readrb -> nios_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_result;         // nios_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_b;              // nios_custom_instruction_master_multi_xconnect:ci_master0_b -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_c;              // nios_custom_instruction_master_multi_xconnect:ci_master0_c -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_done;           // nios_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // nios_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] nios_custom_instruction_master_multi_xconnect_ci_master0_a;              // nios_custom_instruction_master_multi_xconnect:ci_master0_a -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] nios_custom_instruction_master_multi_xconnect_ci_master0_n;              // nios_custom_instruction_master_multi_xconnect:ci_master0_n -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // nios_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // nios_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_clk;            // nios_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // nios_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_start;          // nios_custom_instruction_master_multi_xconnect:ci_master0_start -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // nios_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readra;         // nios_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_reset;          // nios_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] nios_custom_instruction_master_multi_xconnect_ci_master0_datab;          // nios_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // nios_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         nios_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // nios_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_result; // LCD_Driver_0:result -> nios_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_start;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_start -> LCD_Driver_0:start
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> LCD_Driver_0:dataa
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_done;   // LCD_Driver_0:done -> nios_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // nios_custom_instruction_master_multi_slave_translator0:ci_master_clken -> LCD_Driver_0:clk_en
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_reset -> LCD_Driver_0:reset
	wire  [31:0] nios_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // nios_custom_instruction_master_multi_slave_translator0:ci_master_datab -> LCD_Driver_0:datab
	wire         nios_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // nios_custom_instruction_master_multi_slave_translator0:ci_master_clk -> LCD_Driver_0:clk
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                     // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                       // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_chipselect;                                    // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire         mm_interconnect_0_leds_s1_write;                                         // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                      // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                    // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                      // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                        // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                          // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                           // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                       // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         nios_instruction_master_waitrequest;                                     // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [14:0] nios_instruction_master_address;                                         // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                                            // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire  [31:0] nios_instruction_master_readdata;                                        // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         mm_interconnect_0_nios_jtag_debug_module_waitrequest;                    // nios:jtag_debug_module_waitrequest -> mm_interconnect_0:nios_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_writedata;                      // mm_interconnect_0:nios_jtag_debug_module_writedata -> nios:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios_jtag_debug_module_address;                        // mm_interconnect_0:nios_jtag_debug_module_address -> nios:jtag_debug_module_address
	wire         mm_interconnect_0_nios_jtag_debug_module_write;                          // mm_interconnect_0:nios_jtag_debug_module_write -> nios:jtag_debug_module_write
	wire         mm_interconnect_0_nios_jtag_debug_module_read;                           // mm_interconnect_0:nios_jtag_debug_module_read -> nios:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios_jtag_debug_module_readdata;                       // nios:jtag_debug_module_readdata -> mm_interconnect_0:nios_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios_jtag_debug_module_debugaccess;                    // mm_interconnect_0:nios_jtag_debug_module_debugaccess -> nios:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios_jtag_debug_module_byteenable;                     // mm_interconnect_0:nios_jtag_debug_module_byteenable -> nios:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                                   // mm_interconnect_0:memory_s1_writedata -> memory:writedata
	wire  [10:0] mm_interconnect_0_memory_s1_address;                                     // mm_interconnect_0:memory_s1_address -> memory:address
	wire         mm_interconnect_0_memory_s1_chipselect;                                  // mm_interconnect_0:memory_s1_chipselect -> memory:chipselect
	wire         mm_interconnect_0_memory_s1_clken;                                       // mm_interconnect_0:memory_s1_clken -> memory:clken
	wire         mm_interconnect_0_memory_s1_write;                                       // mm_interconnect_0:memory_s1_write -> memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                                    // memory:readdata -> mm_interconnect_0:memory_s1_readdata
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                                  // mm_interconnect_0:memory_s1_byteenable -> memory:byteenable
	wire         nios_data_master_waitrequest;                                            // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire  [31:0] nios_data_master_writedata;                                              // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [14:0] nios_data_master_address;                                                // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire         nios_data_master_write;                                                  // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire         nios_data_master_read;                                                   // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire  [31:0] nios_data_master_readdata;                                               // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_debugaccess;                                            // nios:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire   [3:0] nios_data_master_byteenable;                                             // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                                    // mm_interconnect_0:buttons_s1_address -> buttons:address
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                                   // buttons:readdata -> mm_interconnect_0:buttons_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_d_irq_irq;                                                          // irq_mapper:sender_irq -> nios:d_irq
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [buttons:reset_n, irq_mapper:reset, jtag:rst_n, leds:reset_n, memory:reset, mm_interconnect_0:nios_reset_n_reset_bridge_in_reset_reset, nios:reset_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [memory:reset_req, nios:reset_req, rst_translator:reset_req_in]

	proj_qsys_nios nios (
		.clk                                   (clk_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (nios_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios_data_master_read),                                //                          .read
		.d_readdata                            (nios_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios_data_master_write),                               //                          .write
		.d_writedata                           (nios_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios_instruction_master_read),                         //                          .read
		.i_readdata                            (nios_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_multi_done                       (nios_custom_instruction_master_done),                  // custom_instruction_master.done
		.E_ci_multi_clk_en                     (nios_custom_instruction_master_clk_en),                //                          .clk_en
		.E_ci_multi_start                      (nios_custom_instruction_master_start),                 //                          .start
		.E_ci_result                           (nios_custom_instruction_master_result),                //                          .result
		.D_ci_a                                (nios_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (nios_custom_instruction_master_clk),                   //                          .clk
		.E_ci_multi_reset                      (nios_custom_instruction_master_reset),                 //                          .reset
		.E_ci_multi_reset_req                  (nios_custom_instruction_master_reset_req)              //                          .reset_req
	);

	proj_qsys_memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)      //       .reset_req
	);

	proj_qsys_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	proj_qsys_buttons buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_external_connection_export)     // external_connection.export
	);

	proj_qsys_leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_external_connection_export)       // external_connection.export
	);

	lcd_driver lcd_driver_0 (
		.dataa  (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.clk    (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //                              .clk
		.clk_en (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //                              .clk_en
		.start  (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //                              .start
		.reset  (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //                              .reset
		.done   (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //                              .done
		.result (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //                              .result
		.datab  (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //                              .datab
		.en     (en_export),                                                               //                   conduit_end.export
		.rw     (rw_export),                                                               //                 conduit_end_1.export
		.rs     (rs_export),                                                               //                 conduit_end_2.export
		.db     (db_export)                                                                //                 conduit_end_3.export
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios_custom_instruction_master_translator (
		.ci_slave_dataa            (nios_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                    //                .ipending
		.ci_slave_estatus          (),                                                                    //                .estatus
		.ci_slave_multi_clk        (nios_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                    //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                    //                .datab
		.comb_ci_master_result     (),                                                                    //                .result
		.comb_ci_master_n          (),                                                                    //                .n
		.comb_ci_master_readra     (),                                                                    //                .readra
		.comb_ci_master_readrb     (),                                                                    //                .readrb
		.comb_ci_master_writerc    (),                                                                    //                .writerc
		.comb_ci_master_a          (),                                                                    //                .a
		.comb_ci_master_b          (),                                                                    //                .b
		.comb_ci_master_c          (),                                                                    //                .c
		.comb_ci_master_ipending   (),                                                                    //                .ipending
		.comb_ci_master_estatus    (),                                                                    //                .estatus
		.multi_ci_master_clk       (nios_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                //     (terminated)
		.ci_slave_multi_result     (),                                                                    //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                         //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                            //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                             //     (terminated)
	);

	proj_qsys_nios_custom_instruction_master_multi_xconnect nios_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (nios_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_clk       (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_n         (),                                                                        // (terminated)
		.ci_master_readra    (),                                                                        // (terminated)
		.ci_master_readrb    (),                                                                        // (terminated)
		.ci_master_writerc   (),                                                                        // (terminated)
		.ci_master_a         (),                                                                        // (terminated)
		.ci_master_b         (),                                                                        // (terminated)
		.ci_master_c         (),                                                                        // (terminated)
		.ci_master_ipending  (),                                                                        // (terminated)
		.ci_master_estatus   (),                                                                        // (terminated)
		.ci_master_reset_req ()                                                                         // (terminated)
	);

	proj_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (clk_clk),                                              //                            clk_clk.clk
		.nios_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // nios_reset_n_reset_bridge_in_reset.reset
		.nios_data_master_address                 (nios_data_master_address),                             //                   nios_data_master.address
		.nios_data_master_waitrequest             (nios_data_master_waitrequest),                         //                                   .waitrequest
		.nios_data_master_byteenable              (nios_data_master_byteenable),                          //                                   .byteenable
		.nios_data_master_read                    (nios_data_master_read),                                //                                   .read
		.nios_data_master_readdata                (nios_data_master_readdata),                            //                                   .readdata
		.nios_data_master_write                   (nios_data_master_write),                               //                                   .write
		.nios_data_master_writedata               (nios_data_master_writedata),                           //                                   .writedata
		.nios_data_master_debugaccess             (nios_data_master_debugaccess),                         //                                   .debugaccess
		.nios_instruction_master_address          (nios_instruction_master_address),                      //            nios_instruction_master.address
		.nios_instruction_master_waitrequest      (nios_instruction_master_waitrequest),                  //                                   .waitrequest
		.nios_instruction_master_read             (nios_instruction_master_read),                         //                                   .read
		.nios_instruction_master_readdata         (nios_instruction_master_readdata),                     //                                   .readdata
		.buttons_s1_address                       (mm_interconnect_0_buttons_s1_address),                 //                         buttons_s1.address
		.buttons_s1_readdata                      (mm_interconnect_0_buttons_s1_readdata),                //                                   .readdata
		.jtag_avalon_jtag_slave_address           (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //             jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write             (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                   .write
		.jtag_avalon_jtag_slave_read              (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                   .read
		.jtag_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.leds_s1_address                          (mm_interconnect_0_leds_s1_address),                    //                            leds_s1.address
		.leds_s1_write                            (mm_interconnect_0_leds_s1_write),                      //                                   .write
		.leds_s1_readdata                         (mm_interconnect_0_leds_s1_readdata),                   //                                   .readdata
		.leds_s1_writedata                        (mm_interconnect_0_leds_s1_writedata),                  //                                   .writedata
		.leds_s1_chipselect                       (mm_interconnect_0_leds_s1_chipselect),                 //                                   .chipselect
		.memory_s1_address                        (mm_interconnect_0_memory_s1_address),                  //                          memory_s1.address
		.memory_s1_write                          (mm_interconnect_0_memory_s1_write),                    //                                   .write
		.memory_s1_readdata                       (mm_interconnect_0_memory_s1_readdata),                 //                                   .readdata
		.memory_s1_writedata                      (mm_interconnect_0_memory_s1_writedata),                //                                   .writedata
		.memory_s1_byteenable                     (mm_interconnect_0_memory_s1_byteenable),               //                                   .byteenable
		.memory_s1_chipselect                     (mm_interconnect_0_memory_s1_chipselect),               //                                   .chipselect
		.memory_s1_clken                          (mm_interconnect_0_memory_s1_clken),                    //                                   .clken
		.nios_jtag_debug_module_address           (mm_interconnect_0_nios_jtag_debug_module_address),     //             nios_jtag_debug_module.address
		.nios_jtag_debug_module_write             (mm_interconnect_0_nios_jtag_debug_module_write),       //                                   .write
		.nios_jtag_debug_module_read              (mm_interconnect_0_nios_jtag_debug_module_read),        //                                   .read
		.nios_jtag_debug_module_readdata          (mm_interconnect_0_nios_jtag_debug_module_readdata),    //                                   .readdata
		.nios_jtag_debug_module_writedata         (mm_interconnect_0_nios_jtag_debug_module_writedata),   //                                   .writedata
		.nios_jtag_debug_module_byteenable        (mm_interconnect_0_nios_jtag_debug_module_byteenable),  //                                   .byteenable
		.nios_jtag_debug_module_waitrequest       (mm_interconnect_0_nios_jtag_debug_module_waitrequest), //                                   .waitrequest
		.nios_jtag_debug_module_debugaccess       (mm_interconnect_0_nios_jtag_debug_module_debugaccess)  //                                   .debugaccess
	);

	proj_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_jtag_debug_module_reset_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
